magic
tech sky130A
timestamp 1729054991
<< viali >>
rect -81 535 770 552
rect -81 26 770 43
<< metal1 >>
rect -87 552 776 555
rect -87 535 -81 552
rect 770 535 776 552
rect -87 532 776 535
rect -10 274 -5 300
rect 21 274 26 300
rect 55 280 345 294
rect 394 280 684 294
rect 716 273 721 299
rect 747 273 752 299
rect -87 43 776 46
rect -87 26 -81 43
rect 770 26 776 43
rect -87 23 776 26
<< via1 >>
rect -5 274 21 300
rect 721 273 747 299
<< metal2 >>
rect -5 300 21 305
rect 721 299 747 304
rect 21 274 721 299
rect -5 269 21 274
rect 721 268 747 273
use inverter  inverter_0
timestamp 1729050558
transform 1 0 604 0 1 2
box -27 5 184 568
use inverter  inverter_1
timestamp 1729050558
transform 1 0 -72 0 1 3
box -27 5 184 568
use inverter  inverter_2
timestamp 1729050558
transform 1 0 266 0 1 2
box -27 5 184 568
<< labels >>
flabel viali -69 544 -69 544 0 FreeSans 80 0 0 0 VDD
port 0 nsew
flabel viali -71 34 -71 34 0 FreeSans 80 0 0 0 GND
port 1 nsew
flabel via1 8 286 8 286 0 FreeSans 80 0 0 0 OUT
port 2 nsew
<< end >>
